cdnjn
dj
mn
lp
