module tb();


endmodule


