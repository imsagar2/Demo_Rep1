module tb();
endmodule


