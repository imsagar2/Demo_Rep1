cdnjn
dj
dk
